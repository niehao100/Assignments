module InstructionMemory(addr,data);
  input [31:0] addr;
  output [31:0] data;
  reg [31:0] data;

  always @ (*)
    case(addr[31:2])
      30'h0: data <= 32'h3c044000;
      30'h1: data <= 32'h8c880020;
      30'h2: data <= 32'h8c89001c;
      30'h3: data <= 32'h31080008;
      30'h4: data <= 32'h1008fffc;
      30'h5: data <= 32'h8c880020;
      30'h6: data <= 32'h8c8a001c;
      30'h7: data <= 32'h31080008;
      30'h8: data <= 32'h1008fffc;
      30'h9: data <= 32'h21250000;
      30'ha: data <= 32'h21460000;
      30'hb: data <= 32'hac800008;
      30'hc: data <= 32'h00004027;
      30'hd: data <= 32'h20092710;
      30'he: data <= 32'h01094823;
      30'hf: data <= 32'hac890000;
      30'h10: data <= 32'hac880004;
      30'h11: data <= 32'h20080003;
      30'h12: data <= 32'hac880008;
      30'h13: data <= 32'h20a90000;
      30'h14: data <= 32'h20ca0000;
      30'h15: data <= 32'h012a402a;
      30'h16: data <= 32'h15000003;
      30'h17: data <= 32'h214b0000;
      30'h18: data <= 32'h212a0000;
      30'h19: data <= 32'h21690000;
      30'h1a: data <= 32'h112a0003;
      30'h1b: data <= 32'h11200002;
      30'h1c: data <= 32'h01495022;
      30'h1d: data <= 32'h08000054;
      30'h1e: data <= 32'h21420000;
      30'h1f: data <= 32'hac82000c;
      30'h20: data <= 32'hac820018;
      30'h21: data <= 32'h08000004;
      30'h20000000: data <= 32'h03400008; //�쳣
      30'h20000001: data <= 32'h23bdfff4;
      30'h20000002: data <= 32'hafa80000;
      30'h20000003: data <= 32'hafa90004;
      30'h20000004: data <= 32'hafaa0008;
      30'h20000005: data <= 32'h8c810008;
      30'h20000006: data <= 32'h3021fff9;
      30'h20000007: data <= 32'hac810008;
      30'h20000008: data <= 32'h237b0001;
      30'h20000009: data <= 32'h337b0003;
      30'h2000000a: data <= 32'h20080003;
      30'h2000000b: data <= 32'h111b000d;
      30'h2000000c: data <= 32'h2108ffff;
      30'h2000000d: data <= 32'h111b0008;
      30'h2000000e: data <= 32'h2108ffff;
      30'h2000000f: data <= 32'h111b0003;
      30'h20000010: data <= 32'h20c90000;
      30'h20000011: data <= 32'h200a0700;
      30'h20000012: data <= 32'h0800006c;
      30'h20000013: data <= 32'h00064902;
      30'h20000014: data <= 32'h200a0b00;
      30'h20000015: data <= 32'h0800006c;
      30'h20000016: data <= 32'h20a90000;
      30'h20000017: data <= 32'h200a0d00;
      30'h20000018: data <= 32'h0800006c;
      30'h20000019: data <= 32'h00054902;
      30'h2000001a: data <= 32'h200a0e00;
      30'h2000001b: data <= 32'h3129000f;
      30'h2000001c: data <= 32'h2008000f;
      30'h2000001d: data <= 32'h1109003a;
      30'h2000001e: data <= 32'h2108ffff;
      30'h2000001f: data <= 32'h11090036;
      30'h20000020: data <= 32'h2108ffff;
      30'h20000021: data <= 32'h11090032;
      30'h20000022: data <= 32'h2108ffff;
      30'h20000023: data <= 32'h1109002e;
      30'h20000024: data <= 32'h2108ffff;
      30'h20000025: data <= 32'h1109002a;
      30'h20000026: data <= 32'h2108ffff;
      30'h20000027: data <= 32'h11090026;
      30'h20000028: data <= 32'h2108ffff;
      30'h20000029: data <= 32'h11090022;
      30'h2000002a: data <= 32'h2108ffff;
      30'h2000002b: data <= 32'h1109001e;
      30'h2000002c: data <= 32'h2108ffff;
      30'h2000002d: data <= 32'h1109001a;
      30'h2000002e: data <= 32'h2108ffff;
      30'h2000002f: data <= 32'h11090016;
      30'h20000030: data <= 32'h2108ffff;
      30'h20000031: data <= 32'h11090012;
      30'h20000032: data <= 32'h2108ffff;
      30'h20000033: data <= 32'h1109000e;
      30'h20000034: data <= 32'h2108ffff;
      30'h20000035: data <= 32'h1109000a;
      30'h20000036: data <= 32'h2108ffff;
      30'h20000037: data <= 32'h11090006;
      30'h20000038: data <= 32'h2108ffff;
      30'h20000039: data <= 32'h11090002;
      30'h2000003a: data <= 32'h214800c0;
      30'h2000003b: data <= 32'h08000164;
      30'h2000003c: data <= 32'h214800f9;
      30'h2000003d: data <= 32'h08000164;
      30'h2000003e: data <= 32'h214800a4;
      30'h2000003f: data <= 32'h08000164;
      30'h20000040: data <= 32'h214800b0;
      30'h20000041: data <= 32'h08000164;
      30'h20000042: data <= 32'h21480099;
      30'h20000043: data <= 32'h08000164;
      30'h20000044: data <= 32'h21480092;
      30'h20000045: data <= 32'h08000164;
      30'h20000046: data <= 32'h21480082;
      30'h20000047: data <= 32'h08000164;
      30'h20000048: data <= 32'h214800f8;
      30'h20000049: data <= 32'h08000164;
      30'h2000004a: data <= 32'h21480080;
      30'h2000004b: data <= 32'h08000164;
      30'h2000004c: data <= 32'h21480090;
      30'h2000004d: data <= 32'h08000164;
      30'h2000004e: data <= 32'h21480088;
      30'h2000004f: data <= 32'h08000164;
      30'h20000050: data <= 32'h21480083;
      30'h20000051: data <= 32'h08000164;
      30'h20000052: data <= 32'h214800c6;
      30'h20000053: data <= 32'h08000164;
      30'h20000054: data <= 32'h214800a1;
      30'h20000055: data <= 32'h08000164;
      30'h20000056: data <= 32'h21480086;
      30'h20000057: data <= 32'h08000164;
      30'h20000058: data <= 32'h2148008e;
      30'h20000059: data <= 32'hac880014;
      30'h2000005a: data <= 32'h20080002;
      30'h2000005b: data <= 32'h00280825;
      30'h2000005c: data <= 32'hac810008;
      30'h2000005d: data <= 32'h8fa80000;
      30'h2000005e: data <= 32'h8fa90004;
      30'h2000005f: data <= 32'h8faa0008;
      30'h20000060: data <= 32'h23bd000c;
      30'h20000061: data <= 32'h235afffc;
      30'h20000065: data <= 32'h03400008;
      default: data <= 32'h0;
    endcase
endmodule
