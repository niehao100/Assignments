module KS_ADD(A,B,S,cout,cin);
  input [31:0] A;
  input [31:0] B;
  input cin;
  output [31:0] S;
  output[1:0] cout;
  
  wire [31:0] S;
  wire [1:0] cout;
  
  wire [31:0] P_0,G_0,P_1,G_1,P_2,G_2,P_3,G_3,P_4,G_4,P_5,G_5;
  
  assign P_0[0] = A[0]^B[0]^cin;
  assign G_0[0] = (A[0]|B[0])&cin|(A[0]&B[0])&~cin;
  assign P_0[1] = A[1]^B[1];
  assign G_0[1] = A[1]&B[1];
  assign P_0[2] = A[2]^B[2];
  assign G_0[2] = A[2]&B[2];
  assign P_0[3] = A[3]^B[3];
  assign G_0[3] = A[3]&B[3];
  assign P_0[4] = A[4]^B[4];
  assign G_0[4] = A[4]&B[4];
  assign P_0[5] = A[5]^B[5];
  assign G_0[5] = A[5]&B[5];
  assign P_0[6] = A[6]^B[6];
  assign G_0[6] = A[6]&B[6];
  assign P_0[7] = A[7]^B[7];
  assign G_0[7] = A[7]&B[7];
  assign P_0[8] = A[8]^B[8];
  assign G_0[8] = A[8]&B[8];
  assign P_0[9] = A[9]^B[9];
  assign G_0[9] = A[9]&B[9];
  assign P_0[10] = A[10]^B[10];
  assign G_0[10] = A[10]&B[10];
  assign P_0[11] = A[11]^B[11];
  assign G_0[11] = A[11]&B[11];
  assign P_0[12] = A[12]^B[12];
  assign G_0[12] = A[12]&B[12];
  assign P_0[13] = A[13]^B[13];
  assign G_0[13] = A[13]&B[13];
  assign P_0[14] = A[14]^B[14];
  assign G_0[14] = A[14]&B[14];
  assign P_0[15] = A[15]^B[15];
  assign G_0[15] = A[15]&B[15];
  assign P_0[16] = A[16]^B[16];
  assign G_0[16] = A[16]&B[16];
  assign P_0[17] = A[17]^B[17];
  assign G_0[17] = A[17]&B[17];
  assign P_0[18] = A[18]^B[18];
  assign G_0[18] = A[18]&B[18];
  assign P_0[19] = A[19]^B[19];
  assign G_0[19] = A[19]&B[19];
  assign P_0[20] = A[20]^B[20];
  assign G_0[20] = A[20]&B[20];
  assign P_0[21] = A[21]^B[21];
  assign G_0[21] = A[21]&B[21];
  assign P_0[22] = A[22]^B[22];
  assign G_0[22] = A[22]&B[22];
  assign P_0[23] = A[23]^B[23];
  assign G_0[23] = A[23]&B[23];
  assign P_0[24] = A[24]^B[24];
  assign G_0[24] = A[24]&B[24];
  assign P_0[25] = A[25]^B[25];
  assign G_0[25] = A[25]&B[25];
  assign P_0[26] = A[26]^B[26];
  assign G_0[26] = A[26]&B[26];
  assign P_0[27] = A[27]^B[27];
  assign G_0[27] = A[27]&B[27];
  assign P_0[28] = A[28]^B[28];
  assign G_0[28] = A[28]&B[28];
  assign P_0[29] = A[29]^B[29];
  assign G_0[29] = A[29]&B[29];
  assign P_0[30] = A[30]^B[30];
  assign G_0[30] = A[30]&B[30];
  assign P_0[31] = A[31]^B[31];
  assign G_0[31] = A[31]&B[31];
  
  assign P_1[0] = P_0[0];
  assign G_1[0] = G_0[0];
  assign P_1[1] = P_0[1]&P_0[0];
  assign G_1[1] = (P_0[1]&G_0[0])|G_0[1];
  assign P_1[2] = P_0[2]&P_0[1];
  assign G_1[2] = (P_0[2]&G_0[1])|G_0[2];
  assign P_1[3] = P_0[3]&P_0[2];
  assign G_1[3] = (P_0[3]&G_0[2])|G_0[3];
  assign P_1[4] = P_0[4]&P_0[3];
  assign G_1[4] = (P_0[4]&G_0[3])|G_0[4];
  assign P_1[5] = P_0[5]&P_0[4];
  assign G_1[5] = (P_0[5]&G_0[4])|G_0[5];
  assign P_1[6] = P_0[6]&P_0[5];
  assign G_1[6] = (P_0[6]&G_0[5])|G_0[6];
  assign P_1[7] = P_0[7]&P_0[6];
  assign G_1[7] = (P_0[7]&G_0[6])|G_0[7];
  assign P_1[8] = P_0[8]&P_0[7];
  assign G_1[8] = (P_0[8]&G_0[7])|G_0[8];
  assign P_1[9] = P_0[9]&P_0[8];
  assign G_1[9] = (P_0[9]&G_0[8])|G_0[9];
  assign P_1[10] = P_0[10]&P_0[9];
  assign G_1[10] = (P_0[10]&G_0[9])|G_0[10];
  assign P_1[11] = P_0[11]&P_0[10];
  assign G_1[11] = (P_0[11]&G_0[10])|G_0[11];
  assign P_1[12] = P_0[12]&P_0[11];
  assign G_1[12] = (P_0[12]&G_0[11])|G_0[12];
  assign P_1[13] = P_0[13]&P_0[12];
  assign G_1[13] = (P_0[13]&G_0[12])|G_0[13];
  assign P_1[14] = P_0[14]&P_0[13];
  assign G_1[14] = (P_0[14]&G_0[13])|G_0[14];
  assign P_1[15] = P_0[15]&P_0[14];
  assign G_1[15] = (P_0[15]&G_0[14])|G_0[15];
  assign P_1[16] = P_0[16]&P_0[15];
  assign G_1[16] = (P_0[16]&G_0[15])|G_0[16];
  assign P_1[17] = P_0[17]&P_0[16];
  assign G_1[17] = (P_0[17]&G_0[16])|G_0[17];
  assign P_1[18] = P_0[18]&P_0[17];
  assign G_1[18] = (P_0[18]&G_0[17])|G_0[18];
  assign P_1[19] = P_0[19]&P_0[18];
  assign G_1[19] = (P_0[19]&G_0[18])|G_0[19];
  assign P_1[20] = P_0[20]&P_0[19];
  assign G_1[20] = (P_0[20]&G_0[19])|G_0[20];
  assign P_1[21] = P_0[21]&P_0[20];
  assign G_1[21] = (P_0[21]&G_0[20])|G_0[21];
  assign P_1[22] = P_0[22]&P_0[21];
  assign G_1[22] = (P_0[22]&G_0[21])|G_0[22];
  assign P_1[23] = P_0[23]&P_0[22];
  assign G_1[23] = (P_0[23]&G_0[22])|G_0[23];
  assign P_1[24] = P_0[24]&P_0[23];
  assign G_1[24] = (P_0[24]&G_0[23])|G_0[24];
  assign P_1[25] = P_0[25]&P_0[24];
  assign G_1[25] = (P_0[25]&G_0[24])|G_0[25];
  assign P_1[26] = P_0[26]&P_0[25];
  assign G_1[26] = (P_0[26]&G_0[25])|G_0[26];
  assign P_1[27] = P_0[27]&P_0[26];
  assign G_1[27] = (P_0[27]&G_0[26])|G_0[27];
  assign P_1[28] = P_0[28]&P_0[27];
  assign G_1[28] = (P_0[28]&G_0[27])|G_0[28];
  assign P_1[29] = P_0[29]&P_0[28];
  assign G_1[29] = (P_0[29]&G_0[28])|G_0[29];
  assign P_1[30] = P_0[30]&P_0[29];
  assign G_1[30] = (P_0[30]&G_0[29])|G_0[30];
  assign P_1[31] = P_0[31]&P_0[30];
  assign G_1[31] = (P_0[31]&G_0[30])|G_0[31];
  
  assign P_2[0] = P_1[0];
  assign G_2[0] = G_1[0];
  assign P_2[1] = P_1[1];
  assign G_2[1] = G_1[1];
  assign P_2[2] = P_1[2]&P_1[0];
  assign G_2[2] = (P_1[2]&G_1[0])|G_1[2];
  assign P_2[3] = P_1[3]&P_1[1];
  assign G_2[3] = (P_1[3]&G_1[1])|G_1[3];
  assign P_2[4] = P_1[4]&P_1[2];
  assign G_2[4] = (P_1[4]&G_1[2])|G_1[4];
  assign P_2[5] = P_1[5]&P_1[3];
  assign G_2[5] = (P_1[5]&G_1[3])|G_1[5];
  assign P_2[6] = P_1[6]&P_1[4];
  assign G_2[6] = (P_1[6]&G_1[4])|G_1[6];
  assign P_2[7] = P_1[7]&P_1[5];
  assign G_2[7] = (P_1[7]&G_1[5])|G_1[7];
  assign P_2[8] = P_1[8]&P_1[6];
  assign G_2[8] = (P_1[8]&G_1[6])|G_1[8];
  assign P_2[9] = P_1[9]&P_1[7];
  assign G_2[9] = (P_1[9]&G_1[7])|G_1[9];
  assign P_2[10] = P_1[10]&P_1[8];
  assign G_2[10] = (P_1[10]&G_1[8])|G_1[10];
  assign P_2[11] = P_1[11]&P_1[9];
  assign G_2[11] = (P_1[11]&G_1[9])|G_1[11];
  assign P_2[12] = P_1[12]&P_1[10];
  assign G_2[12] = (P_1[12]&G_1[10])|G_1[12];
  assign P_2[13] = P_1[13]&P_1[11];
  assign G_2[13] = (P_1[13]&G_1[11])|G_1[13];
  assign P_2[14] = P_1[14]&P_1[12];
  assign G_2[14] = (P_1[14]&G_1[12])|G_1[14];
  assign P_2[15] = P_1[15]&P_1[13];
  assign G_2[15] = (P_1[15]&G_1[13])|G_1[15];
  assign P_2[16] = P_1[16]&P_1[14];
  assign G_2[16] = (P_1[16]&G_1[14])|G_1[16];
  assign P_2[17] = P_1[17]&P_1[15];
  assign G_2[17] = (P_1[17]&G_1[15])|G_1[17];
  assign P_2[18] = P_1[18]&P_1[16];
  assign G_2[18] = (P_1[18]&G_1[16])|G_1[18];
  assign P_2[19] = P_1[19]&P_1[17];
  assign G_2[19] = (P_1[19]&G_1[17])|G_1[19];
  assign P_2[20] = P_1[20]&P_1[18];
  assign G_2[20] = (P_1[20]&G_1[18])|G_1[20];
  assign P_2[21] = P_1[21]&P_1[19];
  assign G_2[21] = (P_1[21]&G_1[19])|G_1[21];
  assign P_2[22] = P_1[22]&P_1[20];
  assign G_2[22] = (P_1[22]&G_1[20])|G_1[22];
  assign P_2[23] = P_1[23]&P_1[21];
  assign G_2[23] = (P_1[23]&G_1[21])|G_1[23];
  assign P_2[24] = P_1[24]&P_1[22];
  assign G_2[24] = (P_1[24]&G_1[22])|G_1[24];
  assign P_2[25] = P_1[25]&P_1[23];
  assign G_2[25] = (P_1[25]&G_1[23])|G_1[25];
  assign P_2[26] = P_1[26]&P_1[24];
  assign G_2[26] = (P_1[26]&G_1[24])|G_1[26];
  assign P_2[27] = P_1[27]&P_1[25];
  assign G_2[27] = (P_1[27]&G_1[25])|G_1[27];
  assign P_2[28] = P_1[28]&P_1[26];
  assign G_2[28] = (P_1[28]&G_1[26])|G_1[28];
  assign P_2[29] = P_1[29]&P_1[27];
  assign G_2[29] = (P_1[29]&G_1[27])|G_1[29];
  assign P_2[30] = P_1[30]&P_1[28];
  assign G_2[30] = (P_1[30]&G_1[28])|G_1[30];
  assign P_2[31] = P_1[31]&P_1[29];
  assign G_2[31] = (P_1[31]&G_1[29])|G_1[31];
  
  assign P_3[0] = P_2[0];
  assign G_3[0] = G_2[0];
  assign P_3[1] = P_2[1];
  assign G_3[1] = G_2[1];
  assign P_3[2] = P_2[2];
  assign G_3[2] = G_2[2];
  assign P_3[3] = P_2[3];
  assign G_3[3] = G_2[3];
  assign P_3[4] = P_2[4]&P_2[0];
  assign G_3[4] = (P_2[4]&G_2[0])|G_2[4];
  assign P_3[5] = P_2[5]&P_2[1];
  assign G_3[5] = (P_2[5]&G_2[1])|G_2[5];
  assign P_3[6] = P_2[6]&P_2[2];
  assign G_3[6] = (P_2[6]&G_2[2])|G_2[6];
  assign P_3[7] = P_2[7]&P_2[3];
  assign G_3[7] = (P_2[7]&G_2[3])|G_2[7];
  assign P_3[8] = P_2[8]&P_2[4];
  assign G_3[8] = (P_2[8]&G_2[4])|G_2[8];
  assign P_3[9] = P_2[9]&P_2[5];
  assign G_3[9] = (P_2[9]&G_2[5])|G_2[9];
  assign P_3[10] = P_2[10]&P_2[6];
  assign G_3[10] = (P_2[10]&G_2[6])|G_2[10];
  assign P_3[11] = P_2[11]&P_2[7];
  assign G_3[11] = (P_2[11]&G_2[7])|G_2[11];
  assign P_3[12] = P_2[12]&P_2[8];
  assign G_3[12] = (P_2[12]&G_2[8])|G_2[12];
  assign P_3[13] = P_2[13]&P_2[9];
  assign G_3[13] = (P_2[13]&G_2[9])|G_2[13];
  assign P_3[14] = P_2[14]&P_2[10];
  assign G_3[14] = (P_2[14]&G_2[10])|G_2[14];
  assign P_3[15] = P_2[15]&P_2[11];
  assign G_3[15] = (P_2[15]&G_2[11])|G_2[15];
  assign P_3[16] = P_2[16]&P_2[12];
  assign G_3[16] = (P_2[16]&G_2[12])|G_2[16];
  assign P_3[17] = P_2[17]&P_2[13];
  assign G_3[17] = (P_2[17]&G_2[13])|G_2[17];
  assign P_3[18] = P_2[18]&P_2[14];
  assign G_3[18] = (P_2[18]&G_2[14])|G_2[18];
  assign P_3[19] = P_2[19]&P_2[15];
  assign G_3[19] = (P_2[19]&G_2[15])|G_2[19];
  assign P_3[20] = P_2[20]&P_2[16];
  assign G_3[20] = (P_2[20]&G_2[16])|G_2[20];
  assign P_3[21] = P_2[21]&P_2[17];
  assign G_3[21] = (P_2[21]&G_2[17])|G_2[21];
  assign P_3[22] = P_2[22]&P_2[18];
  assign G_3[22] = (P_2[22]&G_2[18])|G_2[22];
  assign P_3[23] = P_2[23]&P_2[19];
  assign G_3[23] = (P_2[23]&G_2[19])|G_2[23];
  assign P_3[24] = P_2[24]&P_2[20];
  assign G_3[24] = (P_2[24]&G_2[20])|G_2[24];
  assign P_3[25] = P_2[25]&P_2[21];
  assign G_3[25] = (P_2[25]&G_2[21])|G_2[25];
  assign P_3[26] = P_2[26]&P_2[22];
  assign G_3[26] = (P_2[26]&G_2[22])|G_2[26];
  assign P_3[27] = P_2[27]&P_2[23];
  assign G_3[27] = (P_2[27]&G_2[23])|G_2[27];
  assign P_3[28] = P_2[28]&P_2[24];
  assign G_3[28] = (P_2[28]&G_2[24])|G_2[28];
  assign P_3[29] = P_2[29]&P_2[25];
  assign G_3[29] = (P_2[29]&G_2[25])|G_2[29];
  assign P_3[30] = P_2[30]&P_2[26];
  assign G_3[30] = (P_2[30]&G_2[26])|G_2[30];
  assign P_3[31] = P_2[31]&P_2[27];
  assign G_3[31] = (P_2[31]&G_2[27])|G_2[31];
  
  assign P_4[0] = P_3[0];
  assign G_4[0] = G_3[0];
  assign P_4[1] = P_3[1];
  assign G_4[1] = G_3[1];
  assign P_4[2] = P_3[2];
  assign G_4[2] = G_3[2];
  assign P_4[3] = P_3[3];
  assign G_4[3] = G_3[3];
  assign P_4[4] = P_3[4];
  assign G_4[4] = G_3[4];
  assign P_4[5] = P_3[5];
  assign G_4[5] = G_3[5];
  assign P_4[6] = P_3[6];
  assign G_4[6] = G_3[6];
  assign P_4[7] = P_3[7];
  assign G_4[7] = G_3[7];
  assign P_4[8] = P_3[8]&P_3[0];
  assign G_4[8] = (P_3[8]&G_3[0])|G_3[8];
  assign P_4[9] = P_3[9]&P_3[1];
  assign G_4[9] = (P_3[9]&G_3[1])|G_3[9];
  assign P_4[10] = P_3[10]&P_3[2];
  assign G_4[10] = (P_3[10]&G_3[2])|G_3[10];
  assign P_4[11] = P_3[11]&P_3[3];
  assign G_4[11] = (P_3[11]&G_3[3])|G_3[11];
  assign P_4[12] = P_3[12]&P_3[4];
  assign G_4[12] = (P_3[12]&G_3[4])|G_3[12];
  assign P_4[13] = P_3[13]&P_3[5];
  assign G_4[13] = (P_3[13]&G_3[5])|G_3[13];
  assign P_4[14] = P_3[14]&P_3[6];
  assign G_4[14] = (P_3[14]&G_3[6])|G_3[14];
  assign P_4[15] = P_3[15]&P_3[7];
  assign G_4[15] = (P_3[15]&G_3[7])|G_3[15];
  assign P_4[16] = P_3[16]&P_3[8];
  assign G_4[16] = (P_3[16]&G_3[8])|G_3[16];
  assign P_4[17] = P_3[17]&P_3[9];
  assign G_4[17] = (P_3[17]&G_3[9])|G_3[17];
  assign P_4[18] = P_3[18]&P_3[10];
  assign G_4[18] = (P_3[18]&G_3[10])|G_3[18];
  assign P_4[19] = P_3[19]&P_3[11];
  assign G_4[19] = (P_3[19]&G_3[11])|G_3[19];
  assign P_4[20] = P_3[20]&P_3[12];
  assign G_4[20] = (P_3[20]&G_3[12])|G_3[20];
  assign P_4[21] = P_3[21]&P_3[13];
  assign G_4[21] = (P_3[21]&G_3[13])|G_3[21];
  assign P_4[22] = P_3[22]&P_3[14];
  assign G_4[22] = (P_3[22]&G_3[14])|G_3[22];
  assign P_4[23] = P_3[23]&P_3[15];
  assign G_4[23] = (P_3[23]&G_3[15])|G_3[23];
  assign P_4[24] = P_3[24]&P_3[16];
  assign G_4[24] = (P_3[24]&G_3[16])|G_3[24];
  assign P_4[25] = P_3[25]&P_3[17];
  assign G_4[25] = (P_3[25]&G_3[17])|G_3[25];
  assign P_4[26] = P_3[26]&P_3[18];
  assign G_4[26] = (P_3[26]&G_3[18])|G_3[26];
  assign P_4[27] = P_3[27]&P_3[19];
  assign G_4[27] = (P_3[27]&G_3[19])|G_3[27];
  assign P_4[28] = P_3[28]&P_3[20];
  assign G_4[28] = (P_3[28]&G_3[20])|G_3[28];
  assign P_4[29] = P_3[29]&P_3[21];
  assign G_4[29] = (P_3[29]&G_3[21])|G_3[29];
  assign P_4[30] = P_3[30]&P_3[22];
  assign G_4[30] = (P_3[30]&G_3[22])|G_3[30];
  assign P_4[31] = P_3[31]&P_3[23];
  assign G_4[31] = (P_3[31]&G_3[23])|G_3[31];
  
  assign P_5[0] = P_4[0];
  assign G_5[0] = G_4[0];
  assign P_5[1] = P_4[1];
  assign G_5[1] = G_4[1];
  assign P_5[2] = P_4[2];
  assign G_5[2] = G_4[2];
  assign P_5[3] = P_4[3];
  assign G_5[3] = G_4[3];
  assign P_5[4] = P_4[4];
  assign G_5[4] = G_4[4];
  assign P_5[5] = P_4[5];
  assign G_5[5] = G_4[5];
  assign P_5[6] = P_4[6];
  assign G_5[6] = G_4[6];
  assign P_5[7] = P_4[7];
  assign G_5[7] = G_4[7];
  assign P_5[8] = P_4[8];
  assign G_5[8] = G_4[8];
  assign P_5[9] = P_4[9];
  assign G_5[9] = G_4[9];
  assign P_5[10] = P_4[10];
  assign G_5[10] = G_4[10];
  assign P_5[11] = P_4[11];
  assign G_5[11] = G_4[11];
  assign P_5[12] = P_4[12];
  assign G_5[12] = G_4[12];
  assign P_5[13] = P_4[13];
  assign G_5[13] = G_4[13];
  assign P_5[14] = P_4[14];
  assign G_5[14] = G_4[14];
  assign P_5[15] = P_4[15];
  assign G_5[15] = G_4[15];
  assign P_5[16] = P_4[16]&P_4[0];
  assign G_5[16] = (P_4[16]&G_4[0])|G_4[16];
  assign P_5[17] = P_4[17]&P_4[1];
  assign G_5[17] = (P_4[17]&G_4[1])|G_4[17];
  assign P_5[18] = P_4[18]&P_4[2];
  assign G_5[18] = (P_4[18]&G_4[2])|G_4[18];
  assign P_5[19] = P_4[19]&P_4[3];
  assign G_5[19] = (P_4[19]&G_4[3])|G_4[19];
  assign P_5[20] = P_4[20]&P_4[4];
  assign G_5[20] = (P_4[20]&G_4[4])|G_4[20];
  assign P_5[21] = P_4[21]&P_4[5];
  assign G_5[21] = (P_4[21]&G_4[5])|G_4[21];
  assign P_5[22] = P_4[22]&P_4[6];
  assign G_5[22] = (P_4[22]&G_4[6])|G_4[22];
  assign P_5[23] = P_4[23]&P_4[7];
  assign G_5[23] = (P_4[23]&G_4[7])|G_4[23];
  assign P_5[24] = P_4[24]&P_4[8];
  assign G_5[24] = (P_4[24]&G_4[8])|G_4[24];
  assign P_5[25] = P_4[25]&P_4[9];
  assign G_5[25] = (P_4[25]&G_4[9])|G_4[25];
  assign P_5[26] = P_4[26]&P_4[10];
  assign G_5[26] = (P_4[26]&G_4[10])|G_4[26];
  assign P_5[27] = P_4[27]&P_4[11];
  assign G_5[27] = (P_4[27]&G_4[11])|G_4[27];
  assign P_5[28] = P_4[28]&P_4[12];
  assign G_5[28] = (P_4[28]&G_4[12])|G_4[28];
  assign P_5[29] = P_4[29]&P_4[13];
  assign G_5[29] = (P_4[29]&G_4[13])|G_4[29];
  assign P_5[30] = P_4[30]&P_4[14];
  assign G_5[30] = (P_4[30]&G_4[14])|G_4[30];
  assign P_5[31] = P_4[31]&P_4[15];
  assign G_5[31] = (P_4[31]&G_4[15])|G_4[31];
  
  assign S[0] = P_0[0];
  assign S[1] = P_0[1]^G_5[0];
  assign S[2] = P_0[2]^G_5[1];
  assign S[3] = P_0[3]^G_5[2];
  assign S[4] = P_0[4]^G_5[3];
  assign S[5] = P_0[5]^G_5[4];
  assign S[6] = P_0[6]^G_5[5];
  assign S[7] = P_0[7]^G_5[6];
  assign S[8] = P_0[8]^G_5[7];
  assign S[9] = P_0[9]^G_5[8];
  assign S[10] = P_0[10]^G_5[9];
  assign S[11] = P_0[11]^G_5[10];
  assign S[12] = P_0[12]^G_5[11];
  assign S[13] = P_0[13]^G_5[12];
  assign S[14] = P_0[14]^G_5[13];
  assign S[15] = P_0[15]^G_5[14];
  assign S[16] = P_0[16]^G_5[15];
  assign S[17] = P_0[17]^G_5[16];
  assign S[18] = P_0[18]^G_5[17];
  assign S[19] = P_0[19]^G_5[18];
  assign S[20] = P_0[20]^G_5[19];
  assign S[21] = P_0[21]^G_5[20];
  assign S[22] = P_0[22]^G_5[21];
  assign S[23] = P_0[23]^G_5[22];
  assign S[24] = P_0[24]^G_5[23];
  assign S[25] = P_0[25]^G_5[24];
  assign S[26] = P_0[26]^G_5[25];
  assign S[27] = P_0[27]^G_5[26];
  assign S[28] = P_0[28]^G_5[27];
  assign S[29] = P_0[29]^G_5[28];
  assign S[30] = P_0[30]^G_5[29];
  assign S[31] = P_0[31]^G_5[30];
  assign cout[1] = G_5[31];
  assign cout[0] = G_5[30];
endmodule
